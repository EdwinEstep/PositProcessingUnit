/* ----------------- Posit Processing Unit Testbench  -----------------
* 
*  Author:  Edwin Estep
*  Class:   CPE 527
*  
*  This is a testbench to send simple operands through the PPU and
*  collect the results.
*/

module tb_ppu();


endmodule